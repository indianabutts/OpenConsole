module gpu_wb_stage(
		    );


endmodule // gpu_wb_stage
