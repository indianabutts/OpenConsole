module gpu_pc(
	      );


endmodule // gpu_pc
