module gpu_controller(
		      );
endmodule // gpu_controller
