module gpu_alu(
	       );

endmodule;
   
