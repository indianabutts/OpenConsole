module gpu_decode(
		  );


endmodule // gpu_decode
