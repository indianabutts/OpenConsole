module gpu_if_stage(
	      );


endmodule // gpu_if
