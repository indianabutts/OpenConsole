module gpu_if(
	      );


endmodule // gpu_if
