module gpu_registers
                   (
		    
                    );

   
endmodule;
 
