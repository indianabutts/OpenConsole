module gpu_ex(
	      );

endmodule // gpu_ex
