module gpu_opcodes(
		   );

   
parameter NOP
parameter ADD
parameter ADDI
parameter ADDU
parameter ADDIU
parameter SUB
parameter SUBU
parameter MULT
parameter MULTU
parameter DIV
parameter DIVU 
parameter SRL
parameter SRA
parameter SLL
parameter MFHI
parameter MFLO
parameter MTHI
parameter MTLO
parameter AND
parameter OR
parameter NOR
parameter NAND
parameter XOR
parameter CMP
parameter BEQ
parameter BNE
parameter JR
parameter J


endmodule // gpu_opcodes
