module gpu_ex_stage(
	      );

endmodule // gpu_ex
