module gpu_mem_stage(
		     );

endmodule // gpu_mem_stage
